module larger_shell_gtx_bmb7_kintex
(
`include "larger_shell_gtx_shared.vh"
