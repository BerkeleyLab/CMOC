`define SESQUI
module larger_shell_gtx_qf2pre_kintex
(
`include "larger_shell_gtx_shared.vh"
