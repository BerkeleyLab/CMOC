`define LB_HI 14
