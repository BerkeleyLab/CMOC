// parse_vfile  tests/test_1/main_test.v
// module=beam1 instance=beam gvar=cavity_n gcnt=2
// parse_vfile :tests/test_1/main_test.v tests/test_1/beam1.v
`define AUTOMATIC_beam .phase_step(beam_array_phase_step[cavity_n]),\
	.modulo(beam_array_modulo[cavity_n]),\
	.phase_init(beam_array_phase_init[cavity_n])
// module=station instance=cavity gvar=cavity_n gcnt=2
// parse_vfile :tests/test_1/main_test.v tests/test_1/station.v
// module=cav4_elec instance=cav4_elec gvar=None gcnt=None
// parse_vfile :tests/test_1/main_test.v:tests/test_1//sub_dir//station.v tests/test_1/cav4_elec.v
// module=cav4_freq instance=freq gvar=mode_n gcnt=3
// parse_vfile :tests/test_1/main_test.v:tests/test_1//sub_dir//station.v:tests/test_1//sub_dir//cav4_elec.v tests/test_1/cav4_freq.v
// module=test_array instance=piezo_couple gvar=None gcnt=None
// parse_vfile :tests/test_1/main_test.v:tests/test_1//sub_dir//station.v tests/test_1/test_array.v
// found output address in module test_array, base=k_out
`define AUTOMATIC_cavity .cav4_elec_phase_step(cavity_array_cav4_elec_phase_step[cavity_n]),\
	.cav4_elec_modulo(cavity_array_cav4_elec_modulo[cavity_n]),\
	.cav4_elec_trace_reset_we(cavity_array_cav4_elec_trace_reset_we[cavity_n]),\
	.cav4_elec_freq_0_signed_large_port(cavity_array_cav4_elec_freq_0_signed_large_port[cavity_n]),\
	.cav4_elec_freq_1_signed_large_port(cavity_array_cav4_elec_freq_1_signed_large_port[cavity_n]),\
	.cav4_elec_freq_2_signed_large_port(cavity_array_cav4_elec_freq_2_signed_large_port[cavity_n]),\
	.cav4_elec_freq_0_single_cycle(cavity_array_cav4_elec_freq_0_single_cycle[cavity_n]),\
	.cav4_elec_freq_1_single_cycle(cavity_array_cav4_elec_freq_1_single_cycle[cavity_n]),\
	.cav4_elec_freq_2_single_cycle(cavity_array_cav4_elec_freq_2_single_cycle[cavity_n]),\
	.cav4_elec_freq_0_add_write_enable_test(cavity_array_cav4_elec_freq_0_add_write_enable_test[cavity_n]),\
	.cav4_elec_freq_1_add_write_enable_test(cavity_array_cav4_elec_freq_1_add_write_enable_test[cavity_n]),\
	.cav4_elec_freq_2_add_write_enable_test(cavity_array_cav4_elec_freq_2_add_write_enable_test[cavity_n]),\
	.cav4_elec_freq_0_add_write_enable_test_we(cavity_array_cav4_elec_freq_0_add_write_enable_test_we[cavity_n]),\
	.cav4_elec_freq_1_add_write_enable_test_we(cavity_array_cav4_elec_freq_1_add_write_enable_test_we[cavity_n]),\
	.cav4_elec_freq_2_add_write_enable_test_we(cavity_array_cav4_elec_freq_2_add_write_enable_test_we[cavity_n]),\
	.piezo_couple_k_out(cavity_array_piezo_couple_k_out[cavity_n]),\
	.piezo_couple_k_out_addr(cavity_array_piezo_couple_k_out_addr[cavity_n])
// machine-generated by newad.py
`ifdef LB_DECODE_main_test
`include "addr_map_main_test.vh"
`define AUTOMATIC_decode\
wire we_beam_0_phase_step = clk2x_write&(`ADDR_HIT_beam_0_phase_step);\
reg [11:0] beam_0_phase_step=0; always @(posedge clk2x_clk) if (we_beam_0_phase_step) beam_0_phase_step <= clk2x_data;\
wire we_beam_1_phase_step = clk2x_write&(`ADDR_HIT_beam_1_phase_step);\
reg [11:0] beam_1_phase_step=0; always @(posedge clk2x_clk) if (we_beam_1_phase_step) beam_1_phase_step <= clk2x_data;\
wire we_beam_0_modulo = clk2x_write&(`ADDR_HIT_beam_0_modulo);\
reg [11:0] beam_0_modulo=0; always @(posedge clk2x_clk) if (we_beam_0_modulo) beam_0_modulo <= clk2x_data;\
wire we_beam_1_modulo = clk2x_write&(`ADDR_HIT_beam_1_modulo);\
reg [11:0] beam_1_modulo=0; always @(posedge clk2x_clk) if (we_beam_1_modulo) beam_1_modulo <= clk2x_data;\
wire we_beam_0_phase_init = clk2x_write&(`ADDR_HIT_beam_0_phase_init);\
reg [11:0] beam_0_phase_init=0; always @(posedge clk2x_clk) if (we_beam_0_phase_init) beam_0_phase_init <= clk2x_data;\
wire we_beam_1_phase_init = clk2x_write&(`ADDR_HIT_beam_1_phase_init);\
reg [11:0] beam_1_phase_init=0; always @(posedge clk2x_clk) if (we_beam_1_phase_init) beam_1_phase_init <= clk2x_data;\
wire we_cavity_0_cav4_elec_phase_step = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_phase_step);\
reg [31:0] cavity_0_cav4_elec_phase_step=0; always @(posedge clk2x_clk) if (we_cavity_0_cav4_elec_phase_step) cavity_0_cav4_elec_phase_step <= clk2x_data;\
wire we_cavity_1_cav4_elec_phase_step = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_phase_step);\
reg [31:0] cavity_1_cav4_elec_phase_step=0; always @(posedge clk2x_clk) if (we_cavity_1_cav4_elec_phase_step) cavity_1_cav4_elec_phase_step <= clk2x_data;\
wire we_cavity_0_cav4_elec_modulo = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_modulo);\
reg [11:0] cavity_0_cav4_elec_modulo=0; always @(posedge clk2x_clk) if (we_cavity_0_cav4_elec_modulo) cavity_0_cav4_elec_modulo <= clk2x_data;\
wire we_cavity_1_cav4_elec_modulo = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_modulo);\
reg [11:0] cavity_1_cav4_elec_modulo=0; always @(posedge clk2x_clk) if (we_cavity_1_cav4_elec_modulo) cavity_1_cav4_elec_modulo <= clk2x_data;\
wire we_cavity_0_cav4_elec_trace_reset_we = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_trace_reset_we);\
wire cavity_0_cav4_elec_trace_reset_we = we_cavity_0_cav4_elec_trace_reset_we;\
wire we_cavity_1_cav4_elec_trace_reset_we = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_trace_reset_we);\
wire cavity_1_cav4_elec_trace_reset_we = we_cavity_1_cav4_elec_trace_reset_we;\
wire we_cavity_0_cav4_elec_freq_0_signed_large_port = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_freq_0_signed_large_port);\
reg [27:0] cavity_0_cav4_elec_freq_0_signed_large_port=0; always @(posedge clk2x_clk) if (we_cavity_0_cav4_elec_freq_0_signed_large_port) cavity_0_cav4_elec_freq_0_signed_large_port <= clk2x_data;\
wire we_cavity_1_cav4_elec_freq_0_signed_large_port = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_freq_0_signed_large_port);\
reg [27:0] cavity_1_cav4_elec_freq_0_signed_large_port=0; always @(posedge clk2x_clk) if (we_cavity_1_cav4_elec_freq_0_signed_large_port) cavity_1_cav4_elec_freq_0_signed_large_port <= clk2x_data;\
wire we_cavity_0_cav4_elec_freq_1_signed_large_port = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_freq_1_signed_large_port);\
reg [27:0] cavity_0_cav4_elec_freq_1_signed_large_port=0; always @(posedge clk2x_clk) if (we_cavity_0_cav4_elec_freq_1_signed_large_port) cavity_0_cav4_elec_freq_1_signed_large_port <= clk2x_data;\
wire we_cavity_1_cav4_elec_freq_1_signed_large_port = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_freq_1_signed_large_port);\
reg [27:0] cavity_1_cav4_elec_freq_1_signed_large_port=0; always @(posedge clk2x_clk) if (we_cavity_1_cav4_elec_freq_1_signed_large_port) cavity_1_cav4_elec_freq_1_signed_large_port <= clk2x_data;\
wire we_cavity_0_cav4_elec_freq_2_signed_large_port = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_freq_2_signed_large_port);\
reg [27:0] cavity_0_cav4_elec_freq_2_signed_large_port=0; always @(posedge clk2x_clk) if (we_cavity_0_cav4_elec_freq_2_signed_large_port) cavity_0_cav4_elec_freq_2_signed_large_port <= clk2x_data;\
wire we_cavity_1_cav4_elec_freq_2_signed_large_port = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_freq_2_signed_large_port);\
reg [27:0] cavity_1_cav4_elec_freq_2_signed_large_port=0; always @(posedge clk2x_clk) if (we_cavity_1_cav4_elec_freq_2_signed_large_port) cavity_1_cav4_elec_freq_2_signed_large_port <= clk2x_data;\
wire we_cavity_0_cav4_elec_freq_0_single_cycle = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_freq_0_single_cycle);\
reg [1:0] cavity_0_cav4_elec_freq_0_single_cycle=0; always @(posedge clk2x_clk) cavity_0_cav4_elec_freq_0_single_cycle <= we_cavity_0_cav4_elec_freq_0_single_cycle ? clk2x_data[1:0] : 2'b0;\
wire we_cavity_1_cav4_elec_freq_0_single_cycle = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_freq_0_single_cycle);\
reg [1:0] cavity_1_cav4_elec_freq_0_single_cycle=0; always @(posedge clk2x_clk) cavity_1_cav4_elec_freq_0_single_cycle <= we_cavity_1_cav4_elec_freq_0_single_cycle ? clk2x_data[1:0] : 2'b0;\
wire we_cavity_0_cav4_elec_freq_1_single_cycle = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_freq_1_single_cycle);\
reg [1:0] cavity_0_cav4_elec_freq_1_single_cycle=0; always @(posedge clk2x_clk) cavity_0_cav4_elec_freq_1_single_cycle <= we_cavity_0_cav4_elec_freq_1_single_cycle ? clk2x_data[1:0] : 2'b0;\
wire we_cavity_1_cav4_elec_freq_1_single_cycle = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_freq_1_single_cycle);\
reg [1:0] cavity_1_cav4_elec_freq_1_single_cycle=0; always @(posedge clk2x_clk) cavity_1_cav4_elec_freq_1_single_cycle <= we_cavity_1_cav4_elec_freq_1_single_cycle ? clk2x_data[1:0] : 2'b0;\
wire we_cavity_0_cav4_elec_freq_2_single_cycle = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_freq_2_single_cycle);\
reg [1:0] cavity_0_cav4_elec_freq_2_single_cycle=0; always @(posedge clk2x_clk) cavity_0_cav4_elec_freq_2_single_cycle <= we_cavity_0_cav4_elec_freq_2_single_cycle ? clk2x_data[1:0] : 2'b0;\
wire we_cavity_1_cav4_elec_freq_2_single_cycle = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_freq_2_single_cycle);\
reg [1:0] cavity_1_cav4_elec_freq_2_single_cycle=0; always @(posedge clk2x_clk) cavity_1_cav4_elec_freq_2_single_cycle <= we_cavity_1_cav4_elec_freq_2_single_cycle ? clk2x_data[1:0] : 2'b0;\
wire we_cavity_0_cav4_elec_freq_0_add_write_enable_test = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_freq_0_add_write_enable_test);\
wire cavity_0_cav4_elec_freq_0_add_write_enable_test_we = we_cavity_0_cav4_elec_freq_0_add_write_enable_test;\
reg [31:0] cavity_0_cav4_elec_freq_0_add_write_enable_test=0; always @(posedge clk2x_clk) if (we_cavity_0_cav4_elec_freq_0_add_write_enable_test) cavity_0_cav4_elec_freq_0_add_write_enable_test <= clk2x_data;\
wire we_cavity_1_cav4_elec_freq_0_add_write_enable_test = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_freq_0_add_write_enable_test);\
wire cavity_1_cav4_elec_freq_0_add_write_enable_test_we = we_cavity_1_cav4_elec_freq_0_add_write_enable_test;\
reg [31:0] cavity_1_cav4_elec_freq_0_add_write_enable_test=0; always @(posedge clk2x_clk) if (we_cavity_1_cav4_elec_freq_0_add_write_enable_test) cavity_1_cav4_elec_freq_0_add_write_enable_test <= clk2x_data;\
wire we_cavity_0_cav4_elec_freq_1_add_write_enable_test = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_freq_1_add_write_enable_test);\
wire cavity_0_cav4_elec_freq_1_add_write_enable_test_we = we_cavity_0_cav4_elec_freq_1_add_write_enable_test;\
reg [31:0] cavity_0_cav4_elec_freq_1_add_write_enable_test=0; always @(posedge clk2x_clk) if (we_cavity_0_cav4_elec_freq_1_add_write_enable_test) cavity_0_cav4_elec_freq_1_add_write_enable_test <= clk2x_data;\
wire we_cavity_1_cav4_elec_freq_1_add_write_enable_test = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_freq_1_add_write_enable_test);\
wire cavity_1_cav4_elec_freq_1_add_write_enable_test_we = we_cavity_1_cav4_elec_freq_1_add_write_enable_test;\
reg [31:0] cavity_1_cav4_elec_freq_1_add_write_enable_test=0; always @(posedge clk2x_clk) if (we_cavity_1_cav4_elec_freq_1_add_write_enable_test) cavity_1_cav4_elec_freq_1_add_write_enable_test <= clk2x_data;\
wire we_cavity_0_cav4_elec_freq_2_add_write_enable_test = clk2x_write&(`ADDR_HIT_cavity_0_cav4_elec_freq_2_add_write_enable_test);\
wire cavity_0_cav4_elec_freq_2_add_write_enable_test_we = we_cavity_0_cav4_elec_freq_2_add_write_enable_test;\
reg [31:0] cavity_0_cav4_elec_freq_2_add_write_enable_test=0; always @(posedge clk2x_clk) if (we_cavity_0_cav4_elec_freq_2_add_write_enable_test) cavity_0_cav4_elec_freq_2_add_write_enable_test <= clk2x_data;\
wire we_cavity_1_cav4_elec_freq_2_add_write_enable_test = clk2x_write&(`ADDR_HIT_cavity_1_cav4_elec_freq_2_add_write_enable_test);\
wire cavity_1_cav4_elec_freq_2_add_write_enable_test_we = we_cavity_1_cav4_elec_freq_2_add_write_enable_test;\
reg [31:0] cavity_1_cav4_elec_freq_2_add_write_enable_test=0; always @(posedge clk2x_clk) if (we_cavity_1_cav4_elec_freq_2_add_write_enable_test) cavity_1_cav4_elec_freq_2_add_write_enable_test <= clk2x_data;\
wire [9:0] cavity_0_piezo_couple_k_out_addr;\
wire [17:0] cavity_0_piezo_couple_k_out;\
wire we_cavity_0_piezo_couple_k_out = clk2x_write&(`ADDR_HIT_cavity_0_piezo_couple_k_out);\
dpram #(.aw(10),.dw(18)) dp_cavity_0_piezo_couple_k_out(\
	.clka(clk2x_clk), .addra(clk2x_addr[9:0]), .dina(clk2x_data[17:0]), .wena(we_cavity_0_piezo_couple_k_out),\
	.clkb(clk2x_clk), .addrb(cavity_0_piezo_couple_k_out_addr), .doutb(cavity_0_piezo_couple_k_out));\
wire [9:0] cavity_1_piezo_couple_k_out_addr;\
wire [17:0] cavity_1_piezo_couple_k_out;\
wire we_cavity_1_piezo_couple_k_out = clk2x_write&(`ADDR_HIT_cavity_1_piezo_couple_k_out);\
dpram #(.aw(10),.dw(18)) dp_cavity_1_piezo_couple_k_out(\
	.clka(clk2x_clk), .addra(clk2x_addr[9:0]), .dina(clk2x_data[17:0]), .wena(we_cavity_1_piezo_couple_k_out),\
	.clkb(clk2x_clk), .addrb(cavity_1_piezo_couple_k_out_addr), .doutb(cavity_1_piezo_couple_k_out));\
wire we_adc_mmcm = lb_write&(`ADDR_HIT_adc_mmcm);\
reg [1:0] adc_mmcm=0; always @(posedge lb_clk) adc_mmcm <= we_adc_mmcm ? lb_data[1:0] : 2'b0;\
wire [31:0] mirror_out_0;wire mirror_write_0 = lb_write &(`ADDR_HIT_MIRROR);\
dpram #(.aw(`MIRROR_WIDTH),.dw(32)) mirror_0(\
	.clka(lb_clk), .addra(lb_addr[`MIRROR_WIDTH-1:0]), .dina(lb_data[31:0]), .wena(mirror_write_0),\
	.clkb(lb_clk), .addrb(lb_addr[`MIRROR_WIDTH-1:0]), .doutb(mirror_out_0));\

`else
`define AUTOMATIC_self input  [11:0] beam_0_phase_step,\
input  [11:0] beam_1_phase_step,\
input  [11:0] beam_0_modulo,\
input  [11:0] beam_1_modulo,\
input  [11:0] beam_0_phase_init,\
input  [11:0] beam_1_phase_init,\
input  [31:0] cavity_0_cav4_elec_phase_step,\
input  [31:0] cavity_1_cav4_elec_phase_step,\
input  [11:0] cavity_0_cav4_elec_modulo,\
input  [11:0] cavity_1_cav4_elec_modulo,\
input  [0:0] cavity_0_cav4_elec_trace_reset_we,\
input  [0:0] cavity_1_cav4_elec_trace_reset_we,\
input signed [27:0] cavity_0_cav4_elec_freq_0_signed_large_port,\
input signed [27:0] cavity_1_cav4_elec_freq_0_signed_large_port,\
input signed [27:0] cavity_0_cav4_elec_freq_1_signed_large_port,\
input signed [27:0] cavity_1_cav4_elec_freq_1_signed_large_port,\
input signed [27:0] cavity_0_cav4_elec_freq_2_signed_large_port,\
input signed [27:0] cavity_1_cav4_elec_freq_2_signed_large_port,\
input  [1:0] cavity_0_cav4_elec_freq_0_single_cycle,\
input  [1:0] cavity_1_cav4_elec_freq_0_single_cycle,\
input  [1:0] cavity_0_cav4_elec_freq_1_single_cycle,\
input  [1:0] cavity_1_cav4_elec_freq_1_single_cycle,\
input  [1:0] cavity_0_cav4_elec_freq_2_single_cycle,\
input  [1:0] cavity_1_cav4_elec_freq_2_single_cycle,\
input  [31:0] cavity_0_cav4_elec_freq_0_add_write_enable_test,\
input  [31:0] cavity_1_cav4_elec_freq_0_add_write_enable_test,\
input  [31:0] cavity_0_cav4_elec_freq_1_add_write_enable_test,\
input  [31:0] cavity_1_cav4_elec_freq_1_add_write_enable_test,\
input  [31:0] cavity_0_cav4_elec_freq_2_add_write_enable_test,\
input  [31:0] cavity_1_cav4_elec_freq_2_add_write_enable_test,\
input  [0:0] cavity_0_cav4_elec_freq_0_add_write_enable_test_we,\
input  [0:0] cavity_1_cav4_elec_freq_0_add_write_enable_test_we,\
input  [0:0] cavity_0_cav4_elec_freq_1_add_write_enable_test_we,\
input  [0:0] cavity_1_cav4_elec_freq_1_add_write_enable_test_we,\
input  [0:0] cavity_0_cav4_elec_freq_2_add_write_enable_test_we,\
input  [0:0] cavity_1_cav4_elec_freq_2_add_write_enable_test_we,\
input signed [17:0] cavity_0_piezo_couple_k_out,\
input signed [17:0] cavity_1_piezo_couple_k_out,\
output  [9:0] cavity_0_piezo_couple_k_out_addr,\
output  [9:0] cavity_1_piezo_couple_k_out_addr
`define AUTOMATIC_decode
`endif
`define AUTOMATIC_map wire  [11:0] beam_array_phase_step [0:1]; assign beam_array_phase_step[0] = beam_0_phase_step;\
 assign beam_array_phase_step[1] = beam_1_phase_step;\
 wire  [11:0] beam_array_modulo [0:1]; assign beam_array_modulo[0] = beam_0_modulo;\
 assign beam_array_modulo[1] = beam_1_modulo;\
 wire  [11:0] beam_array_phase_init [0:1]; assign beam_array_phase_init[0] = beam_0_phase_init;\
 assign beam_array_phase_init[1] = beam_1_phase_init;\
 wire  [31:0] cavity_array_cav4_elec_phase_step [0:1]; assign cavity_array_cav4_elec_phase_step[0] = cavity_0_cav4_elec_phase_step;\
 assign cavity_array_cav4_elec_phase_step[1] = cavity_1_cav4_elec_phase_step;\
 wire  [11:0] cavity_array_cav4_elec_modulo [0:1]; assign cavity_array_cav4_elec_modulo[0] = cavity_0_cav4_elec_modulo;\
 assign cavity_array_cav4_elec_modulo[1] = cavity_1_cav4_elec_modulo;\
 wire  [0:0] cavity_array_cav4_elec_trace_reset_we [0:1]; assign cavity_array_cav4_elec_trace_reset_we[0] = cavity_0_cav4_elec_trace_reset_we;\
 assign cavity_array_cav4_elec_trace_reset_we[1] = cavity_1_cav4_elec_trace_reset_we;\
 wire signed [27:0] cavity_array_cav4_elec_freq_0_signed_large_port [0:1]; assign cavity_array_cav4_elec_freq_0_signed_large_port[0] = cavity_0_cav4_elec_freq_0_signed_large_port;\
 assign cavity_array_cav4_elec_freq_0_signed_large_port[1] = cavity_1_cav4_elec_freq_0_signed_large_port;\
 wire signed [27:0] cavity_array_cav4_elec_freq_1_signed_large_port [0:1]; assign cavity_array_cav4_elec_freq_1_signed_large_port[0] = cavity_0_cav4_elec_freq_1_signed_large_port;\
 assign cavity_array_cav4_elec_freq_1_signed_large_port[1] = cavity_1_cav4_elec_freq_1_signed_large_port;\
 wire signed [27:0] cavity_array_cav4_elec_freq_2_signed_large_port [0:1]; assign cavity_array_cav4_elec_freq_2_signed_large_port[0] = cavity_0_cav4_elec_freq_2_signed_large_port;\
 assign cavity_array_cav4_elec_freq_2_signed_large_port[1] = cavity_1_cav4_elec_freq_2_signed_large_port;\
 wire  [1:0] cavity_array_cav4_elec_freq_0_single_cycle [0:1]; assign cavity_array_cav4_elec_freq_0_single_cycle[0] = cavity_0_cav4_elec_freq_0_single_cycle;\
 assign cavity_array_cav4_elec_freq_0_single_cycle[1] = cavity_1_cav4_elec_freq_0_single_cycle;\
 wire  [1:0] cavity_array_cav4_elec_freq_1_single_cycle [0:1]; assign cavity_array_cav4_elec_freq_1_single_cycle[0] = cavity_0_cav4_elec_freq_1_single_cycle;\
 assign cavity_array_cav4_elec_freq_1_single_cycle[1] = cavity_1_cav4_elec_freq_1_single_cycle;\
 wire  [1:0] cavity_array_cav4_elec_freq_2_single_cycle [0:1]; assign cavity_array_cav4_elec_freq_2_single_cycle[0] = cavity_0_cav4_elec_freq_2_single_cycle;\
 assign cavity_array_cav4_elec_freq_2_single_cycle[1] = cavity_1_cav4_elec_freq_2_single_cycle;\
 wire  [31:0] cavity_array_cav4_elec_freq_0_add_write_enable_test [0:1]; assign cavity_array_cav4_elec_freq_0_add_write_enable_test[0] = cavity_0_cav4_elec_freq_0_add_write_enable_test;\
 assign cavity_array_cav4_elec_freq_0_add_write_enable_test[1] = cavity_1_cav4_elec_freq_0_add_write_enable_test;\
 wire  [31:0] cavity_array_cav4_elec_freq_1_add_write_enable_test [0:1]; assign cavity_array_cav4_elec_freq_1_add_write_enable_test[0] = cavity_0_cav4_elec_freq_1_add_write_enable_test;\
 assign cavity_array_cav4_elec_freq_1_add_write_enable_test[1] = cavity_1_cav4_elec_freq_1_add_write_enable_test;\
 wire  [31:0] cavity_array_cav4_elec_freq_2_add_write_enable_test [0:1]; assign cavity_array_cav4_elec_freq_2_add_write_enable_test[0] = cavity_0_cav4_elec_freq_2_add_write_enable_test;\
 assign cavity_array_cav4_elec_freq_2_add_write_enable_test[1] = cavity_1_cav4_elec_freq_2_add_write_enable_test;\
 wire  [0:0] cavity_array_cav4_elec_freq_0_add_write_enable_test_we [0:1]; assign cavity_array_cav4_elec_freq_0_add_write_enable_test_we[0] = cavity_0_cav4_elec_freq_0_add_write_enable_test_we;\
 assign cavity_array_cav4_elec_freq_0_add_write_enable_test_we[1] = cavity_1_cav4_elec_freq_0_add_write_enable_test_we;\
 wire  [0:0] cavity_array_cav4_elec_freq_1_add_write_enable_test_we [0:1]; assign cavity_array_cav4_elec_freq_1_add_write_enable_test_we[0] = cavity_0_cav4_elec_freq_1_add_write_enable_test_we;\
 assign cavity_array_cav4_elec_freq_1_add_write_enable_test_we[1] = cavity_1_cav4_elec_freq_1_add_write_enable_test_we;\
 wire  [0:0] cavity_array_cav4_elec_freq_2_add_write_enable_test_we [0:1]; assign cavity_array_cav4_elec_freq_2_add_write_enable_test_we[0] = cavity_0_cav4_elec_freq_2_add_write_enable_test_we;\
 assign cavity_array_cav4_elec_freq_2_add_write_enable_test_we[1] = cavity_1_cav4_elec_freq_2_add_write_enable_test_we;\
 wire signed [17:0] cavity_array_piezo_couple_k_out [0:1]; assign cavity_array_piezo_couple_k_out[0] = cavity_0_piezo_couple_k_out;\
 assign cavity_array_piezo_couple_k_out[1] = cavity_1_piezo_couple_k_out;\
 wire  [9:0] cavity_array_piezo_couple_k_out_addr [0:1]; assign cavity_0_piezo_couple_k_out_addr = cavity_array_piezo_couple_k_out_addr[0];\
 assign cavity_1_piezo_couple_k_out_addr = cavity_array_piezo_couple_k_out_addr[1];\

